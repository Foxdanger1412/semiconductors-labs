** Profile: "SCHEMATIC1-sim5"  [ E:\study\lab4-ahmed\lab4-ahmed\lab4-ahmed-pspicefiles\schematic1\sim5.sim ] 

** Creating circuit file "sim5.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../lab4-ahmed-pspicefiles/lab4-ahmed.lib" 
* From [PSPICE NETLIST] section of C:\Users\engmo\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC LIN 1000 10Hz 10Ghz
.STEP NPN QbreakN(VA) LIST 20,1000 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
