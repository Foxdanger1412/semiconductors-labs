** Profile: "SCHEMATIC1-stage3"  [ E:\study\solid labs\semiconductors-labs\lab1\Reverse bias p-n Junction-PSpiceFiles\SCHEMATIC1\stage3.sim ] 

** Creating circuit file "stage3.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../reverse bias p-n junction-pspicefiles/reverse bias p-n junction.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.STEP V_V5 LIST -9.5 9.5 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
